`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/01/19 18:48:05
// Design Name: 
// Module Name: tb_iic_mux_3
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_iic_mux_3(

    );
    
iic_mux_3(
.SEL_I  (),//[1:0]
.SDA_0_O(),
.SDA_0_I(),
.SDA_0_T(),
.SCL_0_O(),
.SCL_0_I(),
.SCL_0_T(),
.SDA_1_O(),
.SDA_1_I(),
.SDA_1_T(),
.SCL_1_O(),
.SCL_1_I(),
.SCL_1_T(),
.SDA_2_O(),
.SDA_2_I(),
.SDA_2_T(),
.SCL_2_O(),
.SCL_2_I(),
.SCL_2_T(),
.SDA_O  (),
.SDA_I  (),
.SDA_T  (),
.SCL_O  (),
.SCL_I  (),
.SCL_T  ()

);  
    
    
endmodule
