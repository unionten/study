`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/08/19 14:14:22
// Design Name: 
// Module Name: spilt
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module spilt32(
input   [31:0] in    ,
output         out0  , 
output         out1  , 
output         out2  , 
output         out3  , 
output         out4  , 
output         out5  , 
output         out6  , 
output         out7  , 
output         out8  , 
output         out9  , 
output         out10 , 
output         out11 , 
output         out12 , 
output         out13 , 
output         out14 , 
output         out15 , 
output         out16 , 
output         out17 , 
output         out18 , 
output         out19 , 
output         out20 , 
output         out21 , 
output         out22 , 
output         out23 , 
output         out24 , 
output         out25 , 
output         out26 , 
output         out27 , 
output         out28 , 
output         out29 , 
output         out30 , 
output         out31 


);
    
    
    
assign  out0   = in[0    ];
assign  out1   = in[1    ];
assign  out2   = in[2    ];
assign  out3   = in[3    ];
assign  out4   = in[4    ];
assign  out5   = in[5    ];
assign  out6   = in[6    ];
assign  out7   = in[7    ];
assign  out8   = in[8    ];
assign  out9   = in[9    ];
assign  out10  = in[10   ];
assign  out11  = in[11   ];
assign  out12  = in[12   ];
assign  out13  = in[13   ];
assign  out14  = in[14   ];
assign  out15  = in[15   ];
assign  out16  = in[16   ];
assign  out17  = in[17   ];
assign  out18  = in[18   ];
assign  out19  = in[19   ];
assign  out20  = in[20   ];
assign  out21  = in[21   ];
assign  out22  = in[22   ];
assign  out23  = in[23   ];
assign  out24  = in[24   ];
assign  out25  = in[25   ];
assign  out26  = in[26   ];
assign  out27  = in[27   ];
assign  out28  = in[28   ];
assign  out29  = in[29   ];
assign  out30  = in[30   ];
assign  out31  = in[31   ];
    
    
    
    
    
    
endmodule
