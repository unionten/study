`timescale 1ns / 1ps
`define DELAY_OUTGEN(clk,rst,data_in,data_out,DATA_WIDTH,DLY)                                           generate if(DLY==0)begin  assign data_out = data_in; end  else if(DLY==1)begin  (*keep="true"*)reg [DATA_WIDTH-1:0] a_temp = 0; always@(posedge clk) a_temp <= data_in; assign data_out = a_temp ; end  else begin  (*keep="true"*) reg [DATA_WIDTH-1:0] a_temp [DLY-1:0] ;always@(posedge clk) begin  if(rst)a_temp[DLY-1] <= 0; else   a_temp[DLY-1] <= data_in; end  for(i=0;i<=DLY-2;i=i+1)begin  always@(posedge clk)begin  if(rst)begin  a_temp[i] <= 0; end  else begin  a_temp[i] <= a_temp[i+1]; end  end  end  assign data_out = a_temp[0]; end  endgenerate

//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/11/05 14:46:36
// 
//////////////////////////////////////////////////////////////////////////////////


module mux2_signal(
input   [C_WIDTH-1:0]  I0   ,
input   [C_WIDTH-1:0]  I1  ,
input                  S   ,
output   [C_WIDTH-1:0]  O

    );
parameter C_WIDTH = 8; 
    
    
assign  O = (S==0 )? I0 : I1 ;


    
    
endmodule
