`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/01/12 13:55:17
// Design Name: 
// Module Name: num2strb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 

//////////////////////////////////////////////////////////////////////////////////



module num2strb(
input  [$clog2(C_STRB_BIT_NUM)-1:0]  NUM_I  ,//exp : 0 ~ 31
output [C_STRB_BIT_NUM-1:0]        STRB_O 

);
    
parameter C_STRB_BIT_NUM = 32  ;


genvar i;



generate for(i=0;i<C_STRB_BIT_NUM;i=i+1)begin
//assign STRB_O[i] = NUM_I==0 ? 1 : ( NUM_I > i ? 1 : 0 );

assign STRB_O[i] =   (NUM_I-1) >= i ? 1 : 0 ;


end
endgenerate





endmodule

 



//module num2strb(
//input  [$clog2(C_STRB_BIT_NUM):0]  NUM_I  ,
//output [C_STRB_BIT_NUM-1:0]        STRB_O
//
//);
//    
//parameter C_STRB_BIT_NUM = 32  ;
//    
//reg [C_STRB_BIT_NUM-1:0] strb;
//
//assign STRB_O = strb;
//
//
//always@(*)begin
//    case(NUM_I)
//        0:  strb = 32'b00000000000000000000000000000000; 
//        1:  strb = 32'b00000000000000000000000000000001; 
//        2:  strb = 32'b00000000000000000000000000000011; 
//        3:  strb = 32'b00000000000000000000000000000111; 
//        4:  strb = 32'b00000000000000000000000000001111; 
//        5:  strb = 32'b00000000000000000000000000011111; 
//        6:  strb = 32'b00000000000000000000000000111111; 
//        7:  strb = 32'b00000000000000000000000001111111; 
//        8:  strb = 32'b00000000000000000000000011111111; 
//        9:  strb = 32'b00000000000000000000000111111111; 
//        10: strb = 32'b00000000000000000000001111111111; 
//        11: strb = 32'b00000000000000000000011111111111; 
//        12: strb = 32'b00000000000000000000111111111111; 
//        13: strb = 32'b00000000000000000001111111111111; 
//        14: strb = 32'b00000000000000000011111111111111; 
//        15: strb = 32'b00000000000000000111111111111111; 
//        16: strb = 32'b00000000000000001111111111111111; 
//        17: strb = 32'b00000000000000011111111111111111; 
//        18: strb = 32'b00000000000000111111111111111111; 
//        19: strb = 32'b00000000000001111111111111111111; 
//        20: strb = 32'b00000000000011111111111111111111; 
//        21: strb = 32'b00000000000111111111111111111111; 
//        22: strb = 32'b00000000001111111111111111111111; 
//        23: strb = 32'b00000000011111111111111111111111; 
//        24: strb = 32'b00000000111111111111111111111111; 
//        25: strb = 32'b00000001111111111111111111111111; 
//        26: strb = 32'b00000011111111111111111111111111; 
//        27: strb = 32'b00000111111111111111111111111111; 
//        28: strb = 32'b00001111111111111111111111111111; 
//        29: strb = 32'b00011111111111111111111111111111; 
//        30: strb = 32'b00111111111111111111111111111111; 
//        31: strb = 32'b01111111111111111111111111111111; 
//        32: strb = 32'b11111111111111111111111111111111; 
//        default:strb = 32'b11111111111111111111111111111111;  
//    endcase
//end
//   
//  
//endmodule




